library verilog;
use verilog.vl_types.all;
entity naive_bus is
end naive_bus;
