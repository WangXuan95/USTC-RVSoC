module instr_rom(
    input  logic clk, rst_n,
    naive_bus.slave  bus
);
localparam  INSTR_CNT = 30'd81;
wire [0:INSTR_CNT-1] [31:0] instr_rom_cell = {
    32'h00010537,   // 0x00000000
    32'h40050113,   // 0x00000004
    32'h00050513,   // 0x00000008
    32'h00200293,   // 0x0000000c
    32'h00552023,   // 0x00000010
    32'h00100293,   // 0x00000014
    32'h00552223,   // 0x00000018
    32'h00100293,   // 0x0000001c
    32'h00552423,   // 0x00000020
    32'h00000593,   // 0x00000024
    32'h00800613,   // 0x00000028
    32'h00006f33,   // 0x0000002c
    32'h020000ef,   // 0x00000030
    32'h00030fb7,   // 0x00000034
    32'h0fc06f13,   // 0x00000038
    32'h01ef8023,   // 0x0000003c
    32'h00c003b7,   // 0x00000040
    32'hfff38393,   // 0x00000044
    32'hfe039ee3,   // 0x00000048
    32'hfb5ff06f,   // 0x0000004c
    32'h0ec5d863,   // 0x00000050
    32'h0005e333,   // 0x00000054
    32'h000663b3,   // 0x00000058
    32'h006502b3,   // 0x0000005c
    32'h0002a283,   // 0x00000060
    32'h04735463,   // 0x00000064
    32'h00750e33,   // 0x00000068
    32'h000e2e03,   // 0x0000006c
    32'h00735863,   // 0x00000070
    32'h005e4663,   // 0x00000074
    32'hffc38393,   // 0x00000078
    32'hfedff06f,   // 0x0000007c
    32'h00650eb3,   // 0x00000080
    32'h01cea023,   // 0x00000084
    32'h00650e33,   // 0x00000088
    32'h000e2e03,   // 0x0000008c
    32'h00735863,   // 0x00000090
    32'h01c2c663,   // 0x00000094
    32'h00430313,   // 0x00000098
    32'hfedff06f,   // 0x0000009c
    32'h00750eb3,   // 0x000000a0
    32'h01cea023,   // 0x000000a4
    32'hfbdff06f,   // 0x000000a8
    32'h00650eb3,   // 0x000000ac
    32'h005ea023,   // 0x000000b0
    32'hffc10113,   // 0x000000b4
    32'h00112023,   // 0x000000b8
    32'hffc10113,   // 0x000000bc
    32'h00b12023,   // 0x000000c0
    32'hffc10113,   // 0x000000c4
    32'h00c12023,   // 0x000000c8
    32'hffc10113,   // 0x000000cc
    32'h00612023,   // 0x000000d0
    32'hffc30613,   // 0x000000d4
    32'hf79ff0ef,   // 0x000000d8
    32'h00012303,   // 0x000000dc
    32'h00410113,   // 0x000000e0
    32'h00012603,   // 0x000000e4
    32'h00410113,   // 0x000000e8
    32'h00012583,   // 0x000000ec
    32'h00410113,   // 0x000000f0
    32'h00012083,   // 0x000000f4
    32'h00410113,   // 0x000000f8
    32'hffc10113,   // 0x000000fc
    32'h00112023,   // 0x00000100
    32'hffc10113,   // 0x00000104
    32'h00b12023,   // 0x00000108
    32'hffc10113,   // 0x0000010c
    32'h00c12023,   // 0x00000110
    32'hffc10113,   // 0x00000114
    32'h00612023,   // 0x00000118
    32'h00430593,   // 0x0000011c
    32'h00012303,   // 0x00000120
    32'h00410113,   // 0x00000124
    32'h00012603,   // 0x00000128
    32'h00410113,   // 0x0000012c
    32'h00012583,   // 0x00000130
    32'h00410113,   // 0x00000134
    32'h00012083,   // 0x00000138
    32'h00410113,   // 0x0000013c
    32'h00008067    // 0x00000140
};

logic [29:0] cell_rd_addr;

assign bus.rd_gnt = bus.rd_req;
assign bus.wr_gnt = bus.wr_req;
assign cell_rd_addr = bus.rd_addr[31:2];
always @ (posedge clk or negedge rst_n)
    if(~rst_n)
        bus.rd_data <= 0;
    else begin
        if(bus.rd_req)
            bus.rd_data <= (cell_rd_addr>=INSTR_CNT) ? 0 : instr_rom_cell[cell_rd_addr];
        else
            bus.rd_data <= 0;
        end

endmodule

