library verilog;
use verilog.vl_types.all;
entity soc_top_tb is
end soc_top_tb;
